library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.mypak.all;

entity wrapper_vhdl_tb is
end entity wrapper_vhdl_tb;

architecture structural of wrapper_vhdl_tb is
    signal clk : std_logic := '1';
    signal clk_2 : std_logic := '1';
    signal rst : std_logic := '1';
    signal rst_bar : std_logic := '0';
    signal uart : std_logic := '1';
    signal counter : integer := 0;
    signal txd_data : std_logic_vector(7 downto 0);
    signal tx_empty, tx_notemp, tx_en, tx_idle : std_logic;

    signal char : std_logic_vector(7 downto 0) := "00000000";
    signal en : std_logic := '0';
    component wrapper_tb_fifo
        port(
            clk : in std_logic;
            srst : in std_logic;
            din : in std_logic_vector(7 downto 0);
            wr_en : in std_logic;
            rd_en : in std_logic;
            dout : out std_logic_vector(7 downto 0);
            full : out std_logic;
            empty : out std_logic;
            wr_rst_busy : out std_logic;
            rd_rst_busy : out std_logic 
        );
    end component;

    type diff_pair is array(natural range <>) of std_logic_vector(0 to 1);
    signal fmc1_lpc_clk : diff_pair(0 to 1);
    signal fmc1_lpc_la : diff_pair(0 to 33);
    signal fmc1_lpc_scl : std_logic;
    signal fmc1_lpc_sda : std_logic;
    signal fmc2_lpc_clk : diff_pair(0 to 1);
    signal fmc2_lpc_la : diff_pair(0 to 33);
    signal fmc2_lpc_scl : std_logic;
    signal fmc2_lpc_sda : std_logic;
    signal fmc3_hpc_clk : diff_pair(0 to 1);
    signal fmc3_hpc_la : diff_pair(0 to 33);
    signal fmc3_hpc_scl : std_logic;
    signal fmc3_hpc_sda : std_logic;
begin
    clk <= not clk after 2500 ps;
    clk_2 <= not clk_2 after 2000 ps;

    process(clk_2)
    begin
        if rising_edge(clk_2) then
            if rst = '1' then
                counter <= 0;
            else
                counter <= counter + 1;
            end if;
        end if;
    end process;

    input : entity work.uart_tx port map(
        clk => clk_2,
        rst => rst,
        txd_out => uart,
        din => txd_data,
        dval_in => tx_notemp,
        den_out => tx_en,
        idle_out => tx_idle
    );
    tx_notemp <= not tx_empty;

    fifo : wrapper_tb_fifo port map(
        clk => clk_2,
        srst => rst,
        din => char,
        wr_en => en,
        rd_en => tx_en,
        dout => txd_data,
        full => open,
        empty => tx_empty,
        wr_rst_busy => open,
        rd_rst_busy => open
    );

    rst <= '0' after 50000 ns;
    rst_bar <= not rst;

    process(clk_2)
    begin
        if rising_edge(clk_2) then

            -- COMMAND GENERATION START

            if counter = 102 then
                en <= '1';
                char <= x"3a";
            elsif counter = 103 then
                char <= x"42";
            elsif counter = 104 then
                char <= x"55";
            elsif counter = 105 then
                char <= x"53";
            elsif counter = 106 then
                char <= x"5f";
            elsif counter = 107 then
                char <= x"2e";
            elsif counter = 108 then
                char <= x"52";
            elsif counter = 109 then
                char <= x"4f";
            elsif counter = 110 then
                char <= x"55";
            elsif counter = 111 then
                char <= x"54";
            elsif counter = 112 then
                char <= x"2e";
            elsif counter = 113 then
                char <= x"57";
            elsif counter = 114 then
                char <= x"52";
            elsif counter = 115 then
                char <= x"54";
            elsif counter = 116 then
                char <= x"45";
            elsif counter = 117 then
                char <= x"2e";
            elsif counter = 118 then
                char <= x"41";
            elsif counter = 119 then
                char <= x"44";
            elsif counter = 120 then
                char <= x"44";
            elsif counter = 121 then
                char <= x"52";
            elsif counter = 122 then
                char <= x"2e";
            elsif counter = 123 then
                char <= x"00";
            elsif counter = 124 then
                char <= x"00";
            elsif counter = 125 then
                char <= x"00";
            elsif counter = 126 then
                char <= x"00";
            elsif counter = 127 then
                char <= x"2e";
            elsif counter = 128 then
                char <= x"44";
            elsif counter = 129 then
                char <= x"41";
            elsif counter = 130 then
                char <= x"54";
            elsif counter = 131 then
                char <= x"41";
            elsif counter = 132 then
                char <= x"2e";
            elsif counter = 133 then
                char <= x"4d";
            elsif counter = 134 then
                char <= x"4c";
            elsif counter = 135 then
                char <= x"4b";
            elsif counter = 136 then
                char <= x"4a";
            elsif counter = 137 then
                char <= x"21";
            elsif counter = 138 then
                char <= x"3a";
            elsif counter = 139 then
                char <= x"42";
            elsif counter = 140 then
                char <= x"55";
            elsif counter = 141 then
                char <= x"53";
            elsif counter = 142 then
                char <= x"5f";
            elsif counter = 143 then
                char <= x"2e";
            elsif counter = 144 then
                char <= x"4d";
            elsif counter = 145 then
                char <= x"4d";
            elsif counter = 146 then
                char <= x"57";
            elsif counter = 147 then
                char <= x"52";
            elsif counter = 148 then
                char <= x"2e";
            elsif counter = 149 then
                char <= x"43";
            elsif counter = 150 then
                char <= x"54";
            elsif counter = 151 then
                char <= x"52";
            elsif counter = 152 then
                char <= x"4c";
            elsif counter = 153 then
                char <= x"2e";
            elsif counter = 154 then
                char <= x"52";
            elsif counter = 155 then
                char <= x"53";
            elsif counter = 156 then
                char <= x"54";
            elsif counter = 157 then
                char <= x"52";
            elsif counter = 158 then
                char <= x"21";
            elsif counter = 159 then
                char <= x"3a";
            elsif counter = 160 then
                char <= x"42";
            elsif counter = 161 then
                char <= x"55";
            elsif counter = 162 then
                char <= x"53";
            elsif counter = 163 then
                char <= x"5f";
            elsif counter = 164 then
                char <= x"2e";
            elsif counter = 165 then
                char <= x"4d";
            elsif counter = 166 then
                char <= x"4d";
            elsif counter = 167 then
                char <= x"57";
            elsif counter = 168 then
                char <= x"52";
            elsif counter = 169 then
                char <= x"2e";
            elsif counter = 170 then
                char <= x"43";
            elsif counter = 171 then
                char <= x"54";
            elsif counter = 172 then
                char <= x"52";
            elsif counter = 173 then
                char <= x"4c";
            elsif counter = 174 then
                char <= x"2e";
            elsif counter = 175 then
                char <= x"53";
            elsif counter = 176 then
                char <= x"45";
            elsif counter = 177 then
                char <= x"54";
            elsif counter = 178 then
                char <= x"52";
            elsif counter = 179 then
                char <= x"21";
            elsif counter = 180 then
                char <= x"3a";
            elsif counter = 181 then
                char <= x"42";
            elsif counter = 182 then
                char <= x"55";
            elsif counter = 183 then
                char <= x"53";
            elsif counter = 184 then
                char <= x"5f";
            elsif counter = 185 then
                char <= x"2e";
            elsif counter = 186 then
                char <= x"4d";
            elsif counter = 187 then
                char <= x"4d";
            elsif counter = 188 then
                char <= x"57";
            elsif counter = 189 then
                char <= x"52";
            elsif counter = 190 then
                char <= x"2e";
            elsif counter = 191 then
                char <= x"43";
            elsif counter = 192 then
                char <= x"54";
            elsif counter = 193 then
                char <= x"52";
            elsif counter = 194 then
                char <= x"4c";
            elsif counter = 195 then
                char <= x"2e";
            elsif counter = 196 then
                char <= x"52";
            elsif counter = 197 then
                char <= x"53";
            elsif counter = 198 then
                char <= x"54";
            elsif counter = 199 then
                char <= x"43";
            elsif counter = 200 then
                char <= x"21";
            elsif counter = 201 then
                char <= x"3a";
            elsif counter = 202 then
                char <= x"42";
            elsif counter = 203 then
                char <= x"55";
            elsif counter = 204 then
                char <= x"53";
            elsif counter = 205 then
                char <= x"5f";
            elsif counter = 206 then
                char <= x"2e";
            elsif counter = 207 then
                char <= x"4d";
            elsif counter = 208 then
                char <= x"4d";
            elsif counter = 209 then
                char <= x"57";
            elsif counter = 210 then
                char <= x"52";
            elsif counter = 211 then
                char <= x"2e";
            elsif counter = 212 then
                char <= x"43";
            elsif counter = 213 then
                char <= x"54";
            elsif counter = 214 then
                char <= x"52";
            elsif counter = 215 then
                char <= x"4c";
            elsif counter = 216 then
                char <= x"2e";
            elsif counter = 217 then
                char <= x"53";
            elsif counter = 218 then
                char <= x"45";
            elsif counter = 219 then
                char <= x"54";
            elsif counter = 220 then
                char <= x"43";
            elsif counter = 221 then
                char <= x"21";
            elsif counter = 222 then
                char <= x"3a";
            elsif counter = 223 then
                char <= x"42";
            elsif counter = 224 then
                char <= x"55";
            elsif counter = 225 then
                char <= x"53";
            elsif counter = 226 then
                char <= x"5f";
            elsif counter = 227 then
                char <= x"2e";
            elsif counter = 228 then
                char <= x"4d";
            elsif counter = 229 then
                char <= x"4d";
            elsif counter = 230 then
                char <= x"57";
            elsif counter = 231 then
                char <= x"52";
            elsif counter = 232 then
                char <= x"2e";
            elsif counter = 233 then
                char <= x"4d";
            elsif counter = 234 then
                char <= x"49";
            elsif counter = 235 then
                char <= x"53";
            elsif counter = 236 then
                char <= x"43";
            elsif counter = 237 then
                char <= x"2e";
            elsif counter = 238 then
                char <= x"44";
            elsif counter = 239 then
                char <= x"41";
            elsif counter = 240 then
                char <= x"54";
            elsif counter = 241 then
                char <= x"41";
            elsif counter = 242 then
                char <= x"2e";
            elsif counter = 243 then
                char <= x"00";
            elsif counter = 244 then
                char <= x"00";
            elsif counter = 245 then
                char <= x"00";
            elsif counter = 246 then
                char <= x"01";
            elsif counter = 247 then
                char <= x"21";
            elsif counter = 248 then
                char <= x"3a";
            elsif counter = 249 then
                char <= x"42";
            elsif counter = 250 then
                char <= x"55";
            elsif counter = 251 then
                char <= x"53";
            elsif counter = 252 then
                char <= x"5f";
            elsif counter = 253 then
                char <= x"2e";
            elsif counter = 254 then
                char <= x"4d";
            elsif counter = 255 then
                char <= x"4d";
            elsif counter = 256 then
                char <= x"57";
            elsif counter = 257 then
                char <= x"52";
            elsif counter = 258 then
                char <= x"2e";
            elsif counter = 259 then
                char <= x"4d";
            elsif counter = 260 then
                char <= x"49";
            elsif counter = 261 then
                char <= x"53";
            elsif counter = 262 then
                char <= x"43";
            elsif counter = 263 then
                char <= x"2e";
            elsif counter = 264 then
                char <= x"44";
            elsif counter = 265 then
                char <= x"41";
            elsif counter = 266 then
                char <= x"54";
            elsif counter = 267 then
                char <= x"41";
            elsif counter = 268 then
                char <= x"2e";
            elsif counter = 269 then
                char <= x"01";
            elsif counter = 270 then
                char <= x"00";
            elsif counter = 271 then
                char <= x"00";
            elsif counter = 272 then
                char <= x"01";
            elsif counter = 273 then
                char <= x"21";
            elsif counter = 274 then
                char <= x"3a";
            elsif counter = 275 then
                char <= x"42";
            elsif counter = 276 then
                char <= x"55";
            elsif counter = 277 then
                char <= x"53";
            elsif counter = 278 then
                char <= x"5f";
            elsif counter = 279 then
                char <= x"2e";
            elsif counter = 280 then
                char <= x"4d";
            elsif counter = 281 then
                char <= x"4d";
            elsif counter = 282 then
                char <= x"57";
            elsif counter = 283 then
                char <= x"52";
            elsif counter = 284 then
                char <= x"2e";
            elsif counter = 285 then
                char <= x"57";
            elsif counter = 286 then
                char <= x"52";
            elsif counter = 287 then
                char <= x"54";
            elsif counter = 288 then
                char <= x"45";
            elsif counter = 289 then
                char <= x"2e";
            elsif counter = 290 then
                char <= x"41";
            elsif counter = 291 then
                char <= x"44";
            elsif counter = 292 then
                char <= x"44";
            elsif counter = 293 then
                char <= x"52";
            elsif counter = 294 then
                char <= x"2e";
            elsif counter = 295 then
                char <= x"00";
            elsif counter = 296 then
                char <= x"00";
            elsif counter = 297 then
                char <= x"00";
            elsif counter = 298 then
                char <= x"1f";
            elsif counter = 299 then
                char <= x"2e";
            elsif counter = 300 then
                char <= x"44";
            elsif counter = 301 then
                char <= x"41";
            elsif counter = 302 then
                char <= x"54";
            elsif counter = 303 then
                char <= x"41";
            elsif counter = 304 then
                char <= x"2e";
            elsif counter = 305 then
                char <= x"00";
            elsif counter = 306 then
                char <= x"00";
            elsif counter = 307 then
                char <= x"03";
            elsif counter = 308 then
                char <= x"e8";
            elsif counter = 309 then
                char <= x"21";
            elsif counter = 310 then
                char <= x"3a";
            elsif counter = 311 then
                char <= x"42";
            elsif counter = 312 then
                char <= x"55";
            elsif counter = 313 then
                char <= x"53";
            elsif counter = 314 then
                char <= x"5f";
            elsif counter = 315 then
                char <= x"2e";
            elsif counter = 316 then
                char <= x"4d";
            elsif counter = 317 then
                char <= x"4d";
            elsif counter = 318 then
                char <= x"57";
            elsif counter = 319 then
                char <= x"52";
            elsif counter = 320 then
                char <= x"2e";
            elsif counter = 321 then
                char <= x"57";
            elsif counter = 322 then
                char <= x"52";
            elsif counter = 323 then
                char <= x"54";
            elsif counter = 324 then
                char <= x"45";
            elsif counter = 325 then
                char <= x"2e";
            elsif counter = 326 then
                char <= x"41";
            elsif counter = 327 then
                char <= x"44";
            elsif counter = 328 then
                char <= x"44";
            elsif counter = 329 then
                char <= x"52";
            elsif counter = 330 then
                char <= x"2e";
            elsif counter = 331 then
                char <= x"00";
            elsif counter = 332 then
                char <= x"00";
            elsif counter = 333 then
                char <= x"00";
            elsif counter = 334 then
                char <= x"1e";
            elsif counter = 335 then
                char <= x"2e";
            elsif counter = 336 then
                char <= x"44";
            elsif counter = 337 then
                char <= x"41";
            elsif counter = 338 then
                char <= x"54";
            elsif counter = 339 then
                char <= x"41";
            elsif counter = 340 then
                char <= x"2e";
            elsif counter = 341 then
                char <= x"01";
            elsif counter = 342 then
                char <= x"94";
            elsif counter = 343 then
                char <= x"10";
            elsif counter = 344 then
                char <= x"10";
            elsif counter = 345 then
                char <= x"21";
            elsif counter = 346 then
                char <= x"3a";
            elsif counter = 347 then
                char <= x"42";
            elsif counter = 348 then
                char <= x"55";
            elsif counter = 349 then
                char <= x"53";
            elsif counter = 350 then
                char <= x"5f";
            elsif counter = 351 then
                char <= x"2e";
            elsif counter = 352 then
                char <= x"4d";
            elsif counter = 353 then
                char <= x"4d";
            elsif counter = 354 then
                char <= x"57";
            elsif counter = 355 then
                char <= x"52";
            elsif counter = 356 then
                char <= x"2e";
            elsif counter = 357 then
                char <= x"57";
            elsif counter = 358 then
                char <= x"52";
            elsif counter = 359 then
                char <= x"54";
            elsif counter = 360 then
                char <= x"45";
            elsif counter = 361 then
                char <= x"2e";
            elsif counter = 362 then
                char <= x"41";
            elsif counter = 363 then
                char <= x"44";
            elsif counter = 364 then
                char <= x"44";
            elsif counter = 365 then
                char <= x"52";
            elsif counter = 366 then
                char <= x"2e";
            elsif counter = 367 then
                char <= x"00";
            elsif counter = 368 then
                char <= x"00";
            elsif counter = 369 then
                char <= x"00";
            elsif counter = 370 then
                char <= x"1d";
            elsif counter = 371 then
                char <= x"2e";
            elsif counter = 372 then
                char <= x"44";
            elsif counter = 373 then
                char <= x"41";
            elsif counter = 374 then
                char <= x"54";
            elsif counter = 375 then
                char <= x"41";
            elsif counter = 376 then
                char <= x"2e";
            elsif counter = 377 then
                char <= x"00";
            elsif counter = 378 then
                char <= x"00";
            elsif counter = 379 then
                char <= x"00";
            elsif counter = 380 then
                char <= x"00";
            elsif counter = 381 then
                char <= x"21";
            elsif counter = 382 then
                char <= x"3a";
            elsif counter = 383 then
                char <= x"42";
            elsif counter = 384 then
                char <= x"55";
            elsif counter = 385 then
                char <= x"53";
            elsif counter = 386 then
                char <= x"5f";
            elsif counter = 387 then
                char <= x"2e";
            elsif counter = 388 then
                char <= x"4d";
            elsif counter = 389 then
                char <= x"4d";
            elsif counter = 390 then
                char <= x"57";
            elsif counter = 391 then
                char <= x"52";
            elsif counter = 392 then
                char <= x"2e";
            elsif counter = 393 then
                char <= x"57";
            elsif counter = 394 then
                char <= x"52";
            elsif counter = 395 then
                char <= x"54";
            elsif counter = 396 then
                char <= x"45";
            elsif counter = 397 then
                char <= x"2e";
            elsif counter = 398 then
                char <= x"41";
            elsif counter = 399 then
                char <= x"44";
            elsif counter = 400 then
                char <= x"44";
            elsif counter = 401 then
                char <= x"52";
            elsif counter = 402 then
                char <= x"2e";
            elsif counter = 403 then
                char <= x"00";
            elsif counter = 404 then
                char <= x"00";
            elsif counter = 405 then
                char <= x"00";
            elsif counter = 406 then
                char <= x"1c";
            elsif counter = 407 then
                char <= x"2e";
            elsif counter = 408 then
                char <= x"44";
            elsif counter = 409 then
                char <= x"41";
            elsif counter = 410 then
                char <= x"54";
            elsif counter = 411 then
                char <= x"41";
            elsif counter = 412 then
                char <= x"2e";
            elsif counter = 413 then
                char <= x"ff";
            elsif counter = 414 then
                char <= x"ff";
            elsif counter = 415 then
                char <= x"d8";
            elsif counter = 416 then
                char <= x"f0";
            elsif counter = 417 then
                char <= x"21";
            elsif counter = 418 then
                char <= x"3a";
            elsif counter = 419 then
                char <= x"42";
            elsif counter = 420 then
                char <= x"55";
            elsif counter = 421 then
                char <= x"53";
            elsif counter = 422 then
                char <= x"5f";
            elsif counter = 423 then
                char <= x"2e";
            elsif counter = 424 then
                char <= x"4d";
            elsif counter = 425 then
                char <= x"4d";
            elsif counter = 426 then
                char <= x"57";
            elsif counter = 427 then
                char <= x"52";
            elsif counter = 428 then
                char <= x"2e";
            elsif counter = 429 then
                char <= x"57";
            elsif counter = 430 then
                char <= x"52";
            elsif counter = 431 then
                char <= x"54";
            elsif counter = 432 then
                char <= x"45";
            elsif counter = 433 then
                char <= x"2e";
            elsif counter = 434 then
                char <= x"41";
            elsif counter = 435 then
                char <= x"44";
            elsif counter = 436 then
                char <= x"44";
            elsif counter = 437 then
                char <= x"52";
            elsif counter = 438 then
                char <= x"2e";
            elsif counter = 439 then
                char <= x"00";
            elsif counter = 440 then
                char <= x"00";
            elsif counter = 441 then
                char <= x"00";
            elsif counter = 442 then
                char <= x"1b";
            elsif counter = 443 then
                char <= x"2e";
            elsif counter = 444 then
                char <= x"44";
            elsif counter = 445 then
                char <= x"41";
            elsif counter = 446 then
                char <= x"54";
            elsif counter = 447 then
                char <= x"41";
            elsif counter = 448 then
                char <= x"2e";
            elsif counter = 449 then
                char <= x"ff";
            elsif counter = 450 then
                char <= x"fc";
            elsif counter = 451 then
                char <= x"f2";
            elsif counter = 452 then
                char <= x"c0";
            elsif counter = 453 then
                char <= x"21";
            elsif counter = 454 then
                char <= x"3a";
            elsif counter = 455 then
                char <= x"42";
            elsif counter = 456 then
                char <= x"55";
            elsif counter = 457 then
                char <= x"53";
            elsif counter = 458 then
                char <= x"5f";
            elsif counter = 459 then
                char <= x"2e";
            elsif counter = 460 then
                char <= x"4d";
            elsif counter = 461 then
                char <= x"4d";
            elsif counter = 462 then
                char <= x"57";
            elsif counter = 463 then
                char <= x"52";
            elsif counter = 464 then
                char <= x"2e";
            elsif counter = 465 then
                char <= x"57";
            elsif counter = 466 then
                char <= x"52";
            elsif counter = 467 then
                char <= x"54";
            elsif counter = 468 then
                char <= x"45";
            elsif counter = 469 then
                char <= x"2e";
            elsif counter = 470 then
                char <= x"41";
            elsif counter = 471 then
                char <= x"44";
            elsif counter = 472 then
                char <= x"44";
            elsif counter = 473 then
                char <= x"52";
            elsif counter = 474 then
                char <= x"2e";
            elsif counter = 475 then
                char <= x"00";
            elsif counter = 476 then
                char <= x"00";
            elsif counter = 477 then
                char <= x"00";
            elsif counter = 478 then
                char <= x"1a";
            elsif counter = 479 then
                char <= x"2e";
            elsif counter = 480 then
                char <= x"44";
            elsif counter = 481 then
                char <= x"41";
            elsif counter = 482 then
                char <= x"54";
            elsif counter = 483 then
                char <= x"41";
            elsif counter = 484 then
                char <= x"2e";
            elsif counter = 485 then
                char <= x"09";
            elsif counter = 486 then
                char <= x"f4";
            elsif counter = 487 then
                char <= x"ff";
            elsif counter = 488 then
                char <= x"5c";
            elsif counter = 489 then
                char <= x"21";
            elsif counter = 490 then
                char <= x"3a";
            elsif counter = 491 then
                char <= x"42";
            elsif counter = 492 then
                char <= x"55";
            elsif counter = 493 then
                char <= x"53";
            elsif counter = 494 then
                char <= x"5f";
            elsif counter = 495 then
                char <= x"2e";
            elsif counter = 496 then
                char <= x"4d";
            elsif counter = 497 then
                char <= x"4d";
            elsif counter = 498 then
                char <= x"57";
            elsif counter = 499 then
                char <= x"52";
            elsif counter = 500 then
                char <= x"2e";
            elsif counter = 501 then
                char <= x"57";
            elsif counter = 502 then
                char <= x"52";
            elsif counter = 503 then
                char <= x"54";
            elsif counter = 504 then
                char <= x"45";
            elsif counter = 505 then
                char <= x"2e";
            elsif counter = 506 then
                char <= x"41";
            elsif counter = 507 then
                char <= x"44";
            elsif counter = 508 then
                char <= x"44";
            elsif counter = 509 then
                char <= x"52";
            elsif counter = 510 then
                char <= x"2e";
            elsif counter = 511 then
                char <= x"00";
            elsif counter = 512 then
                char <= x"00";
            elsif counter = 513 then
                char <= x"00";
            elsif counter = 514 then
                char <= x"19";
            elsif counter = 515 then
                char <= x"2e";
            elsif counter = 516 then
                char <= x"44";
            elsif counter = 517 then
                char <= x"41";
            elsif counter = 518 then
                char <= x"54";
            elsif counter = 519 then
                char <= x"41";
            elsif counter = 520 then
                char <= x"2e";
            elsif counter = 521 then
                char <= x"4f";
            elsif counter = 522 then
                char <= x"a1";
            elsif counter = 523 then
                char <= x"06";
            elsif counter = 524 then
                char <= x"00";
            elsif counter = 525 then
                char <= x"21";
            elsif counter = 526 then
                char <= x"3a";
            elsif counter = 527 then
                char <= x"42";
            elsif counter = 528 then
                char <= x"55";
            elsif counter = 529 then
                char <= x"53";
            elsif counter = 530 then
                char <= x"5f";
            elsif counter = 531 then
                char <= x"2e";
            elsif counter = 532 then
                char <= x"4d";
            elsif counter = 533 then
                char <= x"4d";
            elsif counter = 534 then
                char <= x"57";
            elsif counter = 535 then
                char <= x"52";
            elsif counter = 536 then
                char <= x"2e";
            elsif counter = 537 then
                char <= x"57";
            elsif counter = 538 then
                char <= x"52";
            elsif counter = 539 then
                char <= x"54";
            elsif counter = 540 then
                char <= x"45";
            elsif counter = 541 then
                char <= x"2e";
            elsif counter = 542 then
                char <= x"41";
            elsif counter = 543 then
                char <= x"44";
            elsif counter = 544 then
                char <= x"44";
            elsif counter = 545 then
                char <= x"52";
            elsif counter = 546 then
                char <= x"2e";
            elsif counter = 547 then
                char <= x"00";
            elsif counter = 548 then
                char <= x"00";
            elsif counter = 549 then
                char <= x"00";
            elsif counter = 550 then
                char <= x"18";
            elsif counter = 551 then
                char <= x"2e";
            elsif counter = 552 then
                char <= x"44";
            elsif counter = 553 then
                char <= x"41";
            elsif counter = 554 then
                char <= x"54";
            elsif counter = 555 then
                char <= x"41";
            elsif counter = 556 then
                char <= x"2e";
            elsif counter = 557 then
                char <= x"00";
            elsif counter = 558 then
                char <= x"30";
            elsif counter = 559 then
                char <= x"0f";
            elsif counter = 560 then
                char <= x"ed";
            elsif counter = 561 then
                char <= x"21";
            elsif counter = 562 then
                char <= x"3a";
            elsif counter = 563 then
                char <= x"42";
            elsif counter = 564 then
                char <= x"55";
            elsif counter = 565 then
                char <= x"53";
            elsif counter = 566 then
                char <= x"5f";
            elsif counter = 567 then
                char <= x"2e";
            elsif counter = 568 then
                char <= x"4d";
            elsif counter = 569 then
                char <= x"4d";
            elsif counter = 570 then
                char <= x"57";
            elsif counter = 571 then
                char <= x"52";
            elsif counter = 572 then
                char <= x"2e";
            elsif counter = 573 then
                char <= x"57";
            elsif counter = 574 then
                char <= x"52";
            elsif counter = 575 then
                char <= x"54";
            elsif counter = 576 then
                char <= x"45";
            elsif counter = 577 then
                char <= x"2e";
            elsif counter = 578 then
                char <= x"41";
            elsif counter = 579 then
                char <= x"44";
            elsif counter = 580 then
                char <= x"44";
            elsif counter = 581 then
                char <= x"52";
            elsif counter = 582 then
                char <= x"2e";
            elsif counter = 583 then
                char <= x"00";
            elsif counter = 584 then
                char <= x"00";
            elsif counter = 585 then
                char <= x"00";
            elsif counter = 586 then
                char <= x"17";
            elsif counter = 587 then
                char <= x"2e";
            elsif counter = 588 then
                char <= x"44";
            elsif counter = 589 then
                char <= x"41";
            elsif counter = 590 then
                char <= x"54";
            elsif counter = 591 then
                char <= x"41";
            elsif counter = 592 then
                char <= x"2e";
            elsif counter = 593 then
                char <= x"01";
            elsif counter = 594 then
                char <= x"40";
            elsif counter = 595 then
                char <= x"03";
            elsif counter = 596 then
                char <= x"f0";
            elsif counter = 597 then
                char <= x"21";
            elsif counter = 598 then
                char <= x"3a";
            elsif counter = 599 then
                char <= x"42";
            elsif counter = 600 then
                char <= x"55";
            elsif counter = 601 then
                char <= x"53";
            elsif counter = 602 then
                char <= x"5f";
            elsif counter = 603 then
                char <= x"2e";
            elsif counter = 604 then
                char <= x"4d";
            elsif counter = 605 then
                char <= x"4d";
            elsif counter = 606 then
                char <= x"57";
            elsif counter = 607 then
                char <= x"52";
            elsif counter = 608 then
                char <= x"2e";
            elsif counter = 609 then
                char <= x"57";
            elsif counter = 610 then
                char <= x"52";
            elsif counter = 611 then
                char <= x"54";
            elsif counter = 612 then
                char <= x"45";
            elsif counter = 613 then
                char <= x"2e";
            elsif counter = 614 then
                char <= x"41";
            elsif counter = 615 then
                char <= x"44";
            elsif counter = 616 then
                char <= x"44";
            elsif counter = 617 then
                char <= x"52";
            elsif counter = 618 then
                char <= x"2e";
            elsif counter = 619 then
                char <= x"00";
            elsif counter = 620 then
                char <= x"00";
            elsif counter = 621 then
                char <= x"00";
            elsif counter = 622 then
                char <= x"16";
            elsif counter = 623 then
                char <= x"2e";
            elsif counter = 624 then
                char <= x"44";
            elsif counter = 625 then
                char <= x"41";
            elsif counter = 626 then
                char <= x"54";
            elsif counter = 627 then
                char <= x"41";
            elsif counter = 628 then
                char <= x"2e";
            elsif counter = 629 then
                char <= x"12";
            elsif counter = 630 then
                char <= x"00";
            elsif counter = 631 then
                char <= x"06";
            elsif counter = 632 then
                char <= x"00";
            elsif counter = 633 then
                char <= x"21";
            elsif counter = 634 then
                char <= x"3a";
            elsif counter = 635 then
                char <= x"42";
            elsif counter = 636 then
                char <= x"55";
            elsif counter = 637 then
                char <= x"53";
            elsif counter = 638 then
                char <= x"5f";
            elsif counter = 639 then
                char <= x"2e";
            elsif counter = 640 then
                char <= x"4d";
            elsif counter = 641 then
                char <= x"4d";
            elsif counter = 642 then
                char <= x"57";
            elsif counter = 643 then
                char <= x"52";
            elsif counter = 644 then
                char <= x"2e";
            elsif counter = 645 then
                char <= x"57";
            elsif counter = 646 then
                char <= x"52";
            elsif counter = 647 then
                char <= x"54";
            elsif counter = 648 then
                char <= x"45";
            elsif counter = 649 then
                char <= x"2e";
            elsif counter = 650 then
                char <= x"41";
            elsif counter = 651 then
                char <= x"44";
            elsif counter = 652 then
                char <= x"44";
            elsif counter = 653 then
                char <= x"52";
            elsif counter = 654 then
                char <= x"2e";
            elsif counter = 655 then
                char <= x"00";
            elsif counter = 656 then
                char <= x"00";
            elsif counter = 657 then
                char <= x"00";
            elsif counter = 658 then
                char <= x"15";
            elsif counter = 659 then
                char <= x"2e";
            elsif counter = 660 then
                char <= x"44";
            elsif counter = 661 then
                char <= x"41";
            elsif counter = 662 then
                char <= x"54";
            elsif counter = 663 then
                char <= x"41";
            elsif counter = 664 then
                char <= x"2e";
            elsif counter = 665 then
                char <= x"3b";
            elsif counter = 666 then
                char <= x"80";
            elsif counter = 667 then
                char <= x"02";
            elsif counter = 668 then
                char <= x"56";
            elsif counter = 669 then
                char <= x"21";
            elsif counter = 670 then
                char <= x"3a";
            elsif counter = 671 then
                char <= x"42";
            elsif counter = 672 then
                char <= x"55";
            elsif counter = 673 then
                char <= x"53";
            elsif counter = 674 then
                char <= x"5f";
            elsif counter = 675 then
                char <= x"2e";
            elsif counter = 676 then
                char <= x"4d";
            elsif counter = 677 then
                char <= x"4d";
            elsif counter = 678 then
                char <= x"57";
            elsif counter = 679 then
                char <= x"52";
            elsif counter = 680 then
                char <= x"2e";
            elsif counter = 681 then
                char <= x"57";
            elsif counter = 682 then
                char <= x"52";
            elsif counter = 683 then
                char <= x"54";
            elsif counter = 684 then
                char <= x"45";
            elsif counter = 685 then
                char <= x"2e";
            elsif counter = 686 then
                char <= x"41";
            elsif counter = 687 then
                char <= x"44";
            elsif counter = 688 then
                char <= x"44";
            elsif counter = 689 then
                char <= x"52";
            elsif counter = 690 then
                char <= x"2e";
            elsif counter = 691 then
                char <= x"00";
            elsif counter = 692 then
                char <= x"00";
            elsif counter = 693 then
                char <= x"00";
            elsif counter = 694 then
                char <= x"14";
            elsif counter = 695 then
                char <= x"2e";
            elsif counter = 696 then
                char <= x"44";
            elsif counter = 697 then
                char <= x"41";
            elsif counter = 698 then
                char <= x"54";
            elsif counter = 699 then
                char <= x"41";
            elsif counter = 700 then
                char <= x"2e";
            elsif counter = 701 then
                char <= x"00";
            elsif counter = 702 then
                char <= x"14";
            elsif counter = 703 then
                char <= x"39";
            elsif counter = 704 then
                char <= x"2a";
            elsif counter = 705 then
                char <= x"21";
            elsif counter = 706 then
                char <= x"3a";
            elsif counter = 707 then
                char <= x"42";
            elsif counter = 708 then
                char <= x"55";
            elsif counter = 709 then
                char <= x"53";
            elsif counter = 710 then
                char <= x"5f";
            elsif counter = 711 then
                char <= x"2e";
            elsif counter = 712 then
                char <= x"4d";
            elsif counter = 713 then
                char <= x"4d";
            elsif counter = 714 then
                char <= x"57";
            elsif counter = 715 then
                char <= x"52";
            elsif counter = 716 then
                char <= x"2e";
            elsif counter = 717 then
                char <= x"57";
            elsif counter = 718 then
                char <= x"52";
            elsif counter = 719 then
                char <= x"54";
            elsif counter = 720 then
                char <= x"45";
            elsif counter = 721 then
                char <= x"2e";
            elsif counter = 722 then
                char <= x"41";
            elsif counter = 723 then
                char <= x"44";
            elsif counter = 724 then
                char <= x"44";
            elsif counter = 725 then
                char <= x"52";
            elsif counter = 726 then
                char <= x"2e";
            elsif counter = 727 then
                char <= x"00";
            elsif counter = 728 then
                char <= x"00";
            elsif counter = 729 then
                char <= x"00";
            elsif counter = 730 then
                char <= x"13";
            elsif counter = 731 then
                char <= x"2e";
            elsif counter = 732 then
                char <= x"44";
            elsif counter = 733 then
                char <= x"41";
            elsif counter = 734 then
                char <= x"54";
            elsif counter = 735 then
                char <= x"41";
            elsif counter = 736 then
                char <= x"2e";
            elsif counter = 737 then
                char <= x"3a";
            elsif counter = 738 then
                char <= x"4f";
            elsif counter = 739 then
                char <= x"17";
            elsif counter = 740 then
                char <= x"53";
            elsif counter = 741 then
                char <= x"21";
            elsif counter = 742 then
                char <= x"3a";
            elsif counter = 743 then
                char <= x"42";
            elsif counter = 744 then
                char <= x"55";
            elsif counter = 745 then
                char <= x"53";
            elsif counter = 746 then
                char <= x"5f";
            elsif counter = 747 then
                char <= x"2e";
            elsif counter = 748 then
                char <= x"4d";
            elsif counter = 749 then
                char <= x"4d";
            elsif counter = 750 then
                char <= x"57";
            elsif counter = 751 then
                char <= x"52";
            elsif counter = 752 then
                char <= x"2e";
            elsif counter = 753 then
                char <= x"57";
            elsif counter = 754 then
                char <= x"52";
            elsif counter = 755 then
                char <= x"54";
            elsif counter = 756 then
                char <= x"45";
            elsif counter = 757 then
                char <= x"2e";
            elsif counter = 758 then
                char <= x"41";
            elsif counter = 759 then
                char <= x"44";
            elsif counter = 760 then
                char <= x"44";
            elsif counter = 761 then
                char <= x"52";
            elsif counter = 762 then
                char <= x"2e";
            elsif counter = 763 then
                char <= x"00";
            elsif counter = 764 then
                char <= x"00";
            elsif counter = 765 then
                char <= x"00";
            elsif counter = 766 then
                char <= x"12";
            elsif counter = 767 then
                char <= x"2e";
            elsif counter = 768 then
                char <= x"44";
            elsif counter = 769 then
                char <= x"41";
            elsif counter = 770 then
                char <= x"54";
            elsif counter = 771 then
                char <= x"41";
            elsif counter = 772 then
                char <= x"2e";
            elsif counter = 773 then
                char <= x"01";
            elsif counter = 774 then
                char <= x"e8";
            elsif counter = 775 then
                char <= x"1c";
            elsif counter = 776 then
                char <= x"9c";
            elsif counter = 777 then
                char <= x"21";
            elsif counter = 778 then
                char <= x"3a";
            elsif counter = 779 then
                char <= x"42";
            elsif counter = 780 then
                char <= x"55";
            elsif counter = 781 then
                char <= x"53";
            elsif counter = 782 then
                char <= x"5f";
            elsif counter = 783 then
                char <= x"2e";
            elsif counter = 784 then
                char <= x"4d";
            elsif counter = 785 then
                char <= x"4d";
            elsif counter = 786 then
                char <= x"57";
            elsif counter = 787 then
                char <= x"52";
            elsif counter = 788 then
                char <= x"2e";
            elsif counter = 789 then
                char <= x"57";
            elsif counter = 790 then
                char <= x"52";
            elsif counter = 791 then
                char <= x"54";
            elsif counter = 792 then
                char <= x"45";
            elsif counter = 793 then
                char <= x"2e";
            elsif counter = 794 then
                char <= x"41";
            elsif counter = 795 then
                char <= x"44";
            elsif counter = 796 then
                char <= x"44";
            elsif counter = 797 then
                char <= x"52";
            elsif counter = 798 then
                char <= x"2e";
            elsif counter = 799 then
                char <= x"00";
            elsif counter = 800 then
                char <= x"00";
            elsif counter = 801 then
                char <= x"00";
            elsif counter = 802 then
                char <= x"11";
            elsif counter = 803 then
                char <= x"2e";
            elsif counter = 804 then
                char <= x"44";
            elsif counter = 805 then
                char <= x"41";
            elsif counter = 806 then
                char <= x"54";
            elsif counter = 807 then
                char <= x"41";
            elsif counter = 808 then
                char <= x"2e";
            elsif counter = 809 then
                char <= x"1c";
            elsif counter = 810 then
                char <= x"9c";
            elsif counter = 811 then
                char <= x"5d";
            elsif counter = 812 then
                char <= x"dc";
            elsif counter = 813 then
                char <= x"21";
            elsif counter = 814 then
                char <= x"3a";
            elsif counter = 815 then
                char <= x"42";
            elsif counter = 816 then
                char <= x"55";
            elsif counter = 817 then
                char <= x"53";
            elsif counter = 818 then
                char <= x"5f";
            elsif counter = 819 then
                char <= x"2e";
            elsif counter = 820 then
                char <= x"4d";
            elsif counter = 821 then
                char <= x"4d";
            elsif counter = 822 then
                char <= x"57";
            elsif counter = 823 then
                char <= x"52";
            elsif counter = 824 then
                char <= x"2e";
            elsif counter = 825 then
                char <= x"57";
            elsif counter = 826 then
                char <= x"52";
            elsif counter = 827 then
                char <= x"54";
            elsif counter = 828 then
                char <= x"45";
            elsif counter = 829 then
                char <= x"2e";
            elsif counter = 830 then
                char <= x"41";
            elsif counter = 831 then
                char <= x"44";
            elsif counter = 832 then
                char <= x"44";
            elsif counter = 833 then
                char <= x"52";
            elsif counter = 834 then
                char <= x"2e";
            elsif counter = 835 then
                char <= x"00";
            elsif counter = 836 then
                char <= x"00";
            elsif counter = 837 then
                char <= x"00";
            elsif counter = 838 then
                char <= x"10";
            elsif counter = 839 then
                char <= x"2e";
            elsif counter = 840 then
                char <= x"44";
            elsif counter = 841 then
                char <= x"41";
            elsif counter = 842 then
                char <= x"54";
            elsif counter = 843 then
                char <= x"41";
            elsif counter = 844 then
                char <= x"2e";
            elsif counter = 845 then
                char <= x"00";
            elsif counter = 846 then
                char <= x"00";
            elsif counter = 847 then
                char <= x"00";
            elsif counter = 848 then
                char <= x"05";
            elsif counter = 849 then
                char <= x"21";
            elsif counter = 850 then
                char <= x"3a";
            elsif counter = 851 then
                char <= x"42";
            elsif counter = 852 then
                char <= x"55";
            elsif counter = 853 then
                char <= x"53";
            elsif counter = 854 then
                char <= x"5f";
            elsif counter = 855 then
                char <= x"2e";
            elsif counter = 856 then
                char <= x"4d";
            elsif counter = 857 then
                char <= x"4d";
            elsif counter = 858 then
                char <= x"57";
            elsif counter = 859 then
                char <= x"52";
            elsif counter = 860 then
                char <= x"2e";
            elsif counter = 861 then
                char <= x"57";
            elsif counter = 862 then
                char <= x"52";
            elsif counter = 863 then
                char <= x"54";
            elsif counter = 864 then
                char <= x"45";
            elsif counter = 865 then
                char <= x"2e";
            elsif counter = 866 then
                char <= x"41";
            elsif counter = 867 then
                char <= x"44";
            elsif counter = 868 then
                char <= x"44";
            elsif counter = 869 then
                char <= x"52";
            elsif counter = 870 then
                char <= x"2e";
            elsif counter = 871 then
                char <= x"00";
            elsif counter = 872 then
                char <= x"00";
            elsif counter = 873 then
                char <= x"00";
            elsif counter = 874 then
                char <= x"10";
            elsif counter = 875 then
                char <= x"2e";
            elsif counter = 876 then
                char <= x"44";
            elsif counter = 877 then
                char <= x"41";
            elsif counter = 878 then
                char <= x"54";
            elsif counter = 879 then
                char <= x"41";
            elsif counter = 880 then
                char <= x"2e";
            elsif counter = 881 then
                char <= x"00";
            elsif counter = 882 then
                char <= x"00";
            elsif counter = 883 then
                char <= x"00";
            elsif counter = 884 then
                char <= x"07";
            elsif counter = 885 then
                char <= x"21";
            elsif counter = 886 then
                char <= x"3a";
            elsif counter = 887 then
                char <= x"42";
            elsif counter = 888 then
                char <= x"55";
            elsif counter = 889 then
                char <= x"53";
            elsif counter = 890 then
                char <= x"5f";
            elsif counter = 891 then
                char <= x"2e";
            elsif counter = 892 then
                char <= x"4d";
            elsif counter = 893 then
                char <= x"4d";
            elsif counter = 894 then
                char <= x"57";
            elsif counter = 895 then
                char <= x"52";
            elsif counter = 896 then
                char <= x"2e";
            elsif counter = 897 then
                char <= x"57";
            elsif counter = 898 then
                char <= x"52";
            elsif counter = 899 then
                char <= x"54";
            elsif counter = 900 then
                char <= x"45";
            elsif counter = 901 then
                char <= x"2e";
            elsif counter = 902 then
                char <= x"41";
            elsif counter = 903 then
                char <= x"44";
            elsif counter = 904 then
                char <= x"44";
            elsif counter = 905 then
                char <= x"52";
            elsif counter = 906 then
                char <= x"2e";
            elsif counter = 907 then
                char <= x"00";
            elsif counter = 908 then
                char <= x"00";
            elsif counter = 909 then
                char <= x"00";
            elsif counter = 910 then
                char <= x"10";
            elsif counter = 911 then
                char <= x"2e";
            elsif counter = 912 then
                char <= x"44";
            elsif counter = 913 then
                char <= x"41";
            elsif counter = 914 then
                char <= x"54";
            elsif counter = 915 then
                char <= x"41";
            elsif counter = 916 then
                char <= x"2e";
            elsif counter = 917 then
                char <= x"00";
            elsif counter = 918 then
                char <= x"00";
            elsif counter = 919 then
                char <= x"00";
            elsif counter = 920 then
                char <= x"06";
            elsif counter = 921 then
                char <= x"21";
            elsif counter = 922 then
                en <= '0';
            end if;

            -- COMMAND GENERATION END

        end if;
    end process;

    dut : entity work.wrapper port map(
        sys_clk_p => clk,
        sys_clk_n => not clk,
        rst => rst_bar,
        led_1_o => open,
        led_2_o => open,
        led_3_o => open,
        led_4_o => open,
        panel_led_1_o => open,
        panel_led_2_o => open,
        uart_txd_o => open,
        uart_rxd_i => uart,
        
        fmc1_lpc_clk0_p_b => fmc1_lpc_clk(0)(0),
        fmc1_lpc_clk0_n_b => fmc1_lpc_clk(0)(1),
        fmc1_lpc_clk1_p_b => fmc1_lpc_clk(1)(0),
        fmc1_lpc_clk1_n_b => fmc1_lpc_clk(1)(1),
        fmc1_lpc_la00_p_b => fmc1_lpc_la(0)(0),
        fmc1_lpc_la00_n_b => fmc1_lpc_la(0)(1),
        fmc1_lpc_la01_p_b => fmc1_lpc_la(1)(0),
        fmc1_lpc_la01_n_b => fmc1_lpc_la(1)(1),
        fmc1_lpc_la02_p_b => fmc1_lpc_la(2)(0),
        fmc1_lpc_la02_n_b => fmc1_lpc_la(2)(1),
        fmc1_lpc_la03_p_b => fmc1_lpc_la(3)(0),
        fmc1_lpc_la03_n_b => fmc1_lpc_la(3)(1),
        fmc1_lpc_la04_p_b => fmc1_lpc_la(4)(0),
        fmc1_lpc_la04_n_b => fmc1_lpc_la(4)(1),
        fmc1_lpc_la05_p_b => fmc1_lpc_la(5)(0),
        fmc1_lpc_la05_n_b => fmc1_lpc_la(5)(1),
        fmc1_lpc_la06_p_b => fmc1_lpc_la(6)(0),
        fmc1_lpc_la06_n_b => fmc1_lpc_la(6)(1),
        fmc1_lpc_la07_p_b => fmc1_lpc_la(7)(0),
        fmc1_lpc_la07_n_b => fmc1_lpc_la(7)(1),
        fmc1_lpc_la08_p_b => fmc1_lpc_la(8)(0),
        fmc1_lpc_la08_n_b => fmc1_lpc_la(8)(1),
        fmc1_lpc_la09_p_b => fmc1_lpc_la(9)(0),
        fmc1_lpc_la09_n_b => fmc1_lpc_la(9)(1),
        fmc1_lpc_la10_p_b => fmc1_lpc_la(10)(0),
        fmc1_lpc_la10_n_b => fmc1_lpc_la(10)(1),
        fmc1_lpc_la11_p_b => fmc1_lpc_la(11)(0),
        fmc1_lpc_la11_n_b => fmc1_lpc_la(11)(1),
        fmc1_lpc_la12_p_b => fmc1_lpc_la(12)(0),
        fmc1_lpc_la12_n_b => fmc1_lpc_la(12)(1),
        fmc1_lpc_la13_p_b => fmc1_lpc_la(13)(0),
        fmc1_lpc_la13_n_b => fmc1_lpc_la(13)(1),
        fmc1_lpc_la14_p_b => fmc1_lpc_la(14)(0),
        fmc1_lpc_la14_n_b => fmc1_lpc_la(14)(1),
        fmc1_lpc_la15_p_b => fmc1_lpc_la(15)(0),
        fmc1_lpc_la15_n_b => fmc1_lpc_la(15)(1),
        fmc1_lpc_la16_p_b => fmc1_lpc_la(16)(0),
        fmc1_lpc_la16_n_b => fmc1_lpc_la(16)(1),
        fmc1_lpc_la17_p_b => fmc1_lpc_la(17)(0),
        fmc1_lpc_la17_n_b => fmc1_lpc_la(17)(1),
        fmc1_lpc_la18_p_b => fmc1_lpc_la(18)(0),
        fmc1_lpc_la18_n_b => fmc1_lpc_la(18)(1),
        fmc1_lpc_la19_p_b => fmc1_lpc_la(19)(0),
        fmc1_lpc_la19_n_b => fmc1_lpc_la(19)(1),
        fmc1_lpc_la20_p_b => fmc1_lpc_la(20)(0),
        fmc1_lpc_la20_n_b => fmc1_lpc_la(20)(1),
        fmc1_lpc_la21_p_b => fmc1_lpc_la(21)(0),
        fmc1_lpc_la21_n_b => fmc1_lpc_la(21)(1),
        fmc1_lpc_la22_p_b => fmc1_lpc_la(22)(0),
        fmc1_lpc_la22_n_b => fmc1_lpc_la(22)(1),
        fmc1_lpc_la23_p_b => fmc1_lpc_la(23)(0),
        fmc1_lpc_la23_n_b => fmc1_lpc_la(23)(1),
        fmc1_lpc_la24_p_b => fmc1_lpc_la(24)(0),
        fmc1_lpc_la24_n_b => fmc1_lpc_la(24)(1),
        fmc1_lpc_la25_p_b => fmc1_lpc_la(25)(0),
        fmc1_lpc_la25_n_b => fmc1_lpc_la(25)(1),
        fmc1_lpc_la26_p_b => fmc1_lpc_la(26)(0),
        fmc1_lpc_la26_n_b => fmc1_lpc_la(26)(1),
        fmc1_lpc_la27_p_b => fmc1_lpc_la(27)(0),
        fmc1_lpc_la27_n_b => fmc1_lpc_la(27)(1),
        fmc1_lpc_la28_p_b => fmc1_lpc_la(28)(0),
        fmc1_lpc_la28_n_b => fmc1_lpc_la(28)(1),
        fmc1_lpc_la29_p_b => fmc1_lpc_la(29)(0),
        fmc1_lpc_la29_n_b => fmc1_lpc_la(29)(1),
        fmc1_lpc_la30_p_b => fmc1_lpc_la(30)(0),
        fmc1_lpc_la30_n_b => fmc1_lpc_la(30)(1),
        fmc1_lpc_la31_p_b => fmc1_lpc_la(31)(0),
        fmc1_lpc_la31_n_b => fmc1_lpc_la(31)(1),
        fmc1_lpc_la32_p_b => fmc1_lpc_la(32)(0),
        fmc1_lpc_la32_n_b => fmc1_lpc_la(32)(1),
        fmc1_lpc_la33_p_b => fmc1_lpc_la(33)(0),
        fmc1_lpc_la33_n_b => fmc1_lpc_la(33)(1),
        fmc1_lpc_scl_b => fmc1_lpc_scl,
        fmc1_lpc_sda_b => fmc1_lpc_sda,
        
        fmc2_lpc_clk0_p_b => fmc2_lpc_clk(0)(0),
        fmc2_lpc_clk0_n_b => fmc2_lpc_clk(0)(1),
        fmc2_lpc_clk1_p_b => fmc2_lpc_clk(1)(0),
        fmc2_lpc_clk1_n_b => fmc2_lpc_clk(1)(1),
        fmc2_lpc_la00_p_b => fmc2_lpc_la(0)(0),
        fmc2_lpc_la00_n_b => fmc2_lpc_la(0)(1),
        fmc2_lpc_la01_p_b => fmc2_lpc_la(1)(0),
        fmc2_lpc_la01_n_b => fmc2_lpc_la(1)(1),
        fmc2_lpc_la02_p_b => fmc2_lpc_la(2)(0),
        fmc2_lpc_la02_n_b => fmc2_lpc_la(2)(1),
        fmc2_lpc_la03_p_b => fmc2_lpc_la(3)(0),
        fmc2_lpc_la03_n_b => fmc2_lpc_la(3)(1),
        fmc2_lpc_la04_p_b => fmc2_lpc_la(4)(0),
        fmc2_lpc_la04_n_b => fmc2_lpc_la(4)(1),
        fmc2_lpc_la05_p_b => fmc2_lpc_la(5)(0),
        fmc2_lpc_la05_n_b => fmc2_lpc_la(5)(1),
        fmc2_lpc_la06_p_b => fmc2_lpc_la(6)(0),
        fmc2_lpc_la06_n_b => fmc2_lpc_la(6)(1),
        fmc2_lpc_la07_p_b => fmc2_lpc_la(7)(0),
        fmc2_lpc_la07_n_b => fmc2_lpc_la(7)(1),
        fmc2_lpc_la08_p_b => fmc2_lpc_la(8)(0),
        fmc2_lpc_la08_n_b => fmc2_lpc_la(8)(1),
        fmc2_lpc_la09_p_b => fmc2_lpc_la(9)(0),
        fmc2_lpc_la09_n_b => fmc2_lpc_la(9)(1),
        fmc2_lpc_la10_p_b => fmc2_lpc_la(10)(0),
        fmc2_lpc_la10_n_b => fmc2_lpc_la(10)(1),
        fmc2_lpc_la11_p_b => fmc2_lpc_la(11)(0),
        fmc2_lpc_la11_n_b => fmc2_lpc_la(11)(1),
        fmc2_lpc_la12_p_b => fmc2_lpc_la(12)(0),
        fmc2_lpc_la12_n_b => fmc2_lpc_la(12)(1),
        fmc2_lpc_la13_p_b => fmc2_lpc_la(13)(0),
        fmc2_lpc_la13_n_b => fmc2_lpc_la(13)(1),
        fmc2_lpc_la14_p_b => fmc2_lpc_la(14)(0),
        fmc2_lpc_la14_n_b => fmc2_lpc_la(14)(1),
        fmc2_lpc_la15_p_b => fmc2_lpc_la(15)(0),
        fmc2_lpc_la15_n_b => fmc2_lpc_la(15)(1),
        fmc2_lpc_la16_p_b => fmc2_lpc_la(16)(0),
        fmc2_lpc_la16_n_b => fmc2_lpc_la(16)(1),
        fmc2_lpc_la17_p_b => fmc2_lpc_la(17)(0),
        fmc2_lpc_la17_n_b => fmc2_lpc_la(17)(1),
        fmc2_lpc_la18_p_b => fmc2_lpc_la(18)(0),
        fmc2_lpc_la18_n_b => fmc2_lpc_la(18)(1),
        fmc2_lpc_la19_p_b => fmc2_lpc_la(19)(0),
        fmc2_lpc_la19_n_b => fmc2_lpc_la(19)(1),
        fmc2_lpc_la20_p_b => fmc2_lpc_la(20)(0),
        fmc2_lpc_la20_n_b => fmc2_lpc_la(20)(1),
        fmc2_lpc_la21_p_b => fmc2_lpc_la(21)(0),
        fmc2_lpc_la21_n_b => fmc2_lpc_la(21)(1),
        fmc2_lpc_la22_p_b => fmc2_lpc_la(22)(0),
        fmc2_lpc_la22_n_b => fmc2_lpc_la(22)(1),
        fmc2_lpc_la23_p_b => fmc2_lpc_la(23)(0),
        fmc2_lpc_la23_n_b => fmc2_lpc_la(23)(1),
        fmc2_lpc_la24_p_b => fmc2_lpc_la(24)(0),
        fmc2_lpc_la24_n_b => fmc2_lpc_la(24)(1),
        fmc2_lpc_la25_p_b => fmc2_lpc_la(25)(0),
        fmc2_lpc_la25_n_b => fmc2_lpc_la(25)(1),
        fmc2_lpc_la26_p_b => fmc2_lpc_la(26)(0),
        fmc2_lpc_la26_n_b => fmc2_lpc_la(26)(1),
        fmc2_lpc_la27_p_b => fmc2_lpc_la(27)(0),
        fmc2_lpc_la27_n_b => fmc2_lpc_la(27)(1),
        fmc2_lpc_la28_p_b => fmc2_lpc_la(28)(0),
        fmc2_lpc_la28_n_b => fmc2_lpc_la(28)(1),
        fmc2_lpc_la29_p_b => fmc2_lpc_la(29)(0),
        fmc2_lpc_la29_n_b => fmc2_lpc_la(29)(1),
        fmc2_lpc_la30_p_b => fmc2_lpc_la(30)(0),
        fmc2_lpc_la30_n_b => fmc2_lpc_la(30)(1),
        fmc2_lpc_la31_p_b => fmc2_lpc_la(31)(0),
        fmc2_lpc_la31_n_b => fmc2_lpc_la(31)(1),
        fmc2_lpc_la32_p_b => fmc2_lpc_la(32)(0),
        fmc2_lpc_la32_n_b => fmc2_lpc_la(32)(1),
        fmc2_lpc_la33_p_b => fmc2_lpc_la(33)(0),
        fmc2_lpc_la33_n_b => fmc2_lpc_la(33)(1),
        fmc2_lpc_scl_b => fmc2_lpc_scl,
        fmc2_lpc_sda_b => fmc2_lpc_sda,

        fmc3_hpc_clk0_p_b => fmc3_hpc_clk(0)(0),
        fmc3_hpc_clk0_n_b => fmc3_hpc_clk(0)(1),
        fmc3_hpc_clk1_p_b => fmc3_hpc_clk(1)(0),
        fmc3_hpc_clk1_n_b => fmc3_hpc_clk(1)(1),
        fmc3_hpc_la00_p_b => fmc3_hpc_la(0)(0),
        fmc3_hpc_la00_n_b => fmc3_hpc_la(0)(1),
        fmc3_hpc_la01_p_b => fmc3_hpc_la(1)(0),
        fmc3_hpc_la01_n_b => fmc3_hpc_la(1)(1),
        fmc3_hpc_la02_p_b => fmc3_hpc_la(2)(0),
        fmc3_hpc_la02_n_b => fmc3_hpc_la(2)(1),
        fmc3_hpc_la03_p_b => fmc3_hpc_la(3)(0),
        fmc3_hpc_la03_n_b => fmc3_hpc_la(3)(1),
        fmc3_hpc_la04_p_b => fmc3_hpc_la(4)(0),
        fmc3_hpc_la04_n_b => fmc3_hpc_la(4)(1),
        fmc3_hpc_la05_p_b => fmc3_hpc_la(5)(0),
        fmc3_hpc_la05_n_b => fmc3_hpc_la(5)(1),
        fmc3_hpc_la06_p_b => fmc3_hpc_la(6)(0),
        fmc3_hpc_la06_n_b => fmc3_hpc_la(6)(1),
        fmc3_hpc_la07_p_b => fmc3_hpc_la(7)(0),
        fmc3_hpc_la07_n_b => fmc3_hpc_la(7)(1),
        fmc3_hpc_la08_p_b => fmc3_hpc_la(8)(0),
        fmc3_hpc_la08_n_b => fmc3_hpc_la(8)(1),
        fmc3_hpc_la09_p_b => fmc3_hpc_la(9)(0),
        fmc3_hpc_la09_n_b => fmc3_hpc_la(9)(1),
        fmc3_hpc_la10_p_b => fmc3_hpc_la(10)(0),
        fmc3_hpc_la10_n_b => fmc3_hpc_la(10)(1),
        fmc3_hpc_la11_p_b => fmc3_hpc_la(11)(0),
        fmc3_hpc_la11_n_b => fmc3_hpc_la(11)(1),
        fmc3_hpc_la12_p_b => fmc3_hpc_la(12)(0),
        fmc3_hpc_la12_n_b => fmc3_hpc_la(12)(1),
        fmc3_hpc_la13_p_b => fmc3_hpc_la(13)(0),
        fmc3_hpc_la13_n_b => fmc3_hpc_la(13)(1),
        fmc3_hpc_la14_p_b => fmc3_hpc_la(14)(0),
        fmc3_hpc_la14_n_b => fmc3_hpc_la(14)(1),
        fmc3_hpc_la15_p_b => fmc3_hpc_la(15)(0),
        fmc3_hpc_la15_n_b => fmc3_hpc_la(15)(1),
        fmc3_hpc_la16_p_b => fmc3_hpc_la(16)(0),
        fmc3_hpc_la16_n_b => fmc3_hpc_la(16)(1),
        fmc3_hpc_la17_p_b => fmc3_hpc_la(17)(0),
        fmc3_hpc_la17_n_b => fmc3_hpc_la(17)(1),
        fmc3_hpc_la18_p_b => fmc3_hpc_la(18)(0),
        fmc3_hpc_la18_n_b => fmc3_hpc_la(18)(1),
        fmc3_hpc_la19_p_b => fmc3_hpc_la(19)(0),
        fmc3_hpc_la19_n_b => fmc3_hpc_la(19)(1),
        fmc3_hpc_la20_p_b => fmc3_hpc_la(20)(0),
        fmc3_hpc_la20_n_b => fmc3_hpc_la(20)(1),
        fmc3_hpc_la21_p_b => fmc3_hpc_la(21)(0),
        fmc3_hpc_la21_n_b => fmc3_hpc_la(21)(1),
        fmc3_hpc_la22_p_b => fmc3_hpc_la(22)(0),
        fmc3_hpc_la22_n_b => fmc3_hpc_la(22)(1),
        fmc3_hpc_la23_p_b => fmc3_hpc_la(23)(0),
        fmc3_hpc_la23_n_b => fmc3_hpc_la(23)(1),
        fmc3_hpc_la24_p_b => fmc3_hpc_la(24)(0),
        fmc3_hpc_la24_n_b => fmc3_hpc_la(24)(1),
        fmc3_hpc_la25_p_b => fmc3_hpc_la(25)(0),
        fmc3_hpc_la25_n_b => fmc3_hpc_la(25)(1),
        fmc3_hpc_la26_p_b => fmc3_hpc_la(26)(0),
        fmc3_hpc_la26_n_b => fmc3_hpc_la(26)(1),
        fmc3_hpc_la27_p_b => fmc3_hpc_la(27)(0),
        fmc3_hpc_la27_n_b => fmc3_hpc_la(27)(1),
        fmc3_hpc_la28_p_b => fmc3_hpc_la(28)(0),
        fmc3_hpc_la28_n_b => fmc3_hpc_la(28)(1),
        fmc3_hpc_la29_p_b => fmc3_hpc_la(29)(0),
        fmc3_hpc_la29_n_b => fmc3_hpc_la(29)(1),
        fmc3_hpc_la30_p_b => fmc3_hpc_la(30)(0),
        fmc3_hpc_la30_n_b => fmc3_hpc_la(30)(1),
        fmc3_hpc_la31_p_b => fmc3_hpc_la(31)(0),
        fmc3_hpc_la31_n_b => fmc3_hpc_la(31)(1),
        fmc3_hpc_la32_p_b => fmc3_hpc_la(32)(0),
        fmc3_hpc_la32_n_b => fmc3_hpc_la(32)(1),
        fmc3_hpc_la33_p_b => fmc3_hpc_la(33)(0),
        fmc3_hpc_la33_n_b => fmc3_hpc_la(33)(1),
        fmc3_hpc_scl_b => fmc3_hpc_scl,
        fmc3_hpc_sda_b => fmc3_hpc_sda
    );
end architecture structural; 
